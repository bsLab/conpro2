
-- 
-- Definition of  par_FUN_parity3
-- 
--      Fri Dec 19 11:31:38 2008
--      
--      LeonardoSpectrum Level 3, 2005b.24
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity par_FUN_parity3 is
   port (
      REG_RET_FUN_parity3_p_WR : OUT std_logic ;
      REG_RET_FUN_parity3_p_WE : OUT std_logic ;
      REG_ARG_FUN_parity3_x_RD : IN std_logic_vector (63 DOWNTO 0) ;
      PRO_FUN_parity3_ENABLE : IN std_logic ;
      PRO_FUN_parity3_END : OUT std_logic ;
      conpro_system_clk : IN std_logic ;
      conpro_system_reset : IN std_logic) ;
end par_FUN_parity3 ;

architecture main of par_FUN_parity3 is
   signal PRO_FUN_parity3_END_EXMPLR, REG_RET_FUN_parity3_p_WE_EXMPLR, 
      pro_state_66, pro_state_65, pro_state_64, pro_state_63, pro_state_62, 
      pro_state_61, pro_state_60, pro_state_59, pro_state_58, pro_state_57, 
      pro_state_56, pro_state_55, pro_state_54, pro_state_53, pro_state_52, 
      pro_state_51, pro_state_50, pro_state_49, pro_state_48, pro_state_47, 
      pro_state_46, pro_state_45, pro_state_44, pro_state_43, pro_state_42, 
      pro_state_41, pro_state_40, pro_state_39, pro_state_38, pro_state_37, 
      pro_state_36, pro_state_35, pro_state_34, pro_state_33, pro_state_32, 
      pro_state_31, pro_state_30, pro_state_29, pro_state_28, pro_state_27, 
      pro_state_26, pro_state_25, pro_state_24, pro_state_23, pro_state_22, 
      pro_state_21, pro_state_20, pro_state_19, pro_state_18, pro_state_17, 
      pro_state_16, pro_state_15, pro_state_14, pro_state_13, pro_state_12, 
      pro_state_11, pro_state_10, pro_state_9, pro_state_8, pro_state_7, 
      pro_state_6, pro_state_5, pro_state_4, pro_state_3, pro_state_2, 
      pro_state_1, pro_state_0, nx2, nx12, nx22, nx32, nx42, nx52, nx62, 
      nx72, nx82, nx92, nx102, nx112, nx122, nx132, nx142, nx152, nx162, 
      nx172, nx182, nx192, nx202, nx212, nx222, nx232, nx242, nx252, nx262, 
      nx272, nx282, nx292, nx302, nx312, nx322, nx332, nx342, nx352, nx362, 
      nx372, nx382, nx392, nx402, nx412, nx422, nx432, nx442, nx452, nx462, 
      nx472, nx482, nx492, nx502, nx512, nx522, nx532, nx542, nx552, nx562, 
      nx572, nx582, nx592, nx602, nx612, nx622, nx632, nx642, nx652, nx662, 
      nx672, pl, nx684, nx706, xl_0, nx708, nx712, nx720, xl_1, nx726, nx734, 
      xl_2, nx742, nx750, xl_3, nx756, nx764, xl_4, nx774, nx782, xl_5, 
      nx788, nx796, xl_6, nx804, nx812, xl_7, nx818, nx826, xl_8, nx838, 
      nx846, xl_9, nx852, nx860, xl_10, nx868, nx876, xl_11, nx882, nx890, 
      xl_12, nx900, nx908, xl_13, nx914, nx922, xl_14, nx930, nx938, xl_15, 
      nx944, nx952, nx962, xl_16, nx966, nx974, xl_17, nx980, nx988, xl_18, 
      nx996, nx1004, xl_19, nx1010, nx1018, xl_20, nx1028, nx1036, xl_21, 
      nx1042, nx1050, xl_22, nx1058, nx1066, xl_23, nx1072, nx1080, xl_24, 
      nx1092, nx1100, xl_25, nx1106, nx1114, xl_26, nx1122, nx1130, xl_27, 
      nx1136, nx1144, xl_28, nx1154, nx1162, xl_29, nx1168, nx1176, xl_30, 
      nx1184, nx1192, xl_31, nx1198, nx1206, nx1216, xl_32, nx1222, nx1230, 
      xl_33, nx1236, nx1244, xl_34, nx1252, nx1260, xl_35, nx1266, nx1274, 
      xl_36, nx1284, nx1292, xl_37, nx1298, nx1306, xl_38, nx1314, nx1322, 
      xl_39, nx1328, nx1336, xl_40, nx1348, nx1356, xl_41, nx1362, nx1370, 
      xl_42, nx1378, nx1386, xl_43, nx1392, nx1400, xl_44, nx1410, nx1418, 
      xl_45, nx1424, nx1432, xl_46, nx1440, nx1448, xl_47, nx1454, nx1462, 
      nx1472, xl_48, nx1476, nx1484, xl_49, nx1490, nx1498, xl_50, nx1506, 
      nx1514, xl_51, nx1520, nx1528, xl_52, nx1538, nx1546, xl_53, nx1552, 
      nx1560, xl_54, nx1568, nx1576, xl_55, nx1582, nx1590, xl_56, nx1602, 
      nx1610, xl_57, nx1616, nx1624, xl_58, nx1632, nx1640, xl_59, nx1646, 
      nx1654, xl_60, nx1664, nx1672, xl_61, nx1678, nx1686, xl_62, nx1694, 
      nx1702, xl_63, nx1708, nx1716, nx1726, nx1734, nx3346, nx3349, nx3364, 
      nx3378, nx3392, nx3407, nx3421, nx3435, nx3449, nx3464, nx3478, nx3492, 
      nx3506, nx3521, nx3535, nx3549, nx3563, nx3578, nx3582, nx3589, nx3591, 
      nx3593, nx3595, nx3597, nx3599, nx3601, nx3603, nx3605, nx3607, nx3609, 
      nx3611, nx3613, nx3615, nx3617, nx3619, nx3621, nx3623, nx3625, nx3627, 
      nx3629, nx3631, nx3633, nx3635, nx3637, nx3639, nx3641, nx3643, nx3645, 
      nx3647: std_logic ;

begin
   REG_RET_FUN_parity3_p_WE <= REG_RET_FUN_parity3_p_WE_EXMPLR ;
   PRO_FUN_parity3_END <= PRO_FUN_parity3_END_EXMPLR ;
   ix1743 : a2_x2 port map ( q=>REG_RET_FUN_parity3_p_WR, i0=>
      REG_RET_FUN_parity3_p_WE_EXMPLR, i1=>nx3613);
   reg_pro_state_67 : sff1_x4 port map ( q=>REG_RET_FUN_parity3_p_WE_EXMPLR, 
      i=>nx672, ck=>conpro_system_clk);
   reg_pro_state_66 : sff1_x4 port map ( q=>pro_state_66, i=>nx662, ck=>
      conpro_system_clk);
   reg_pro_state_65 : sff1_x4 port map ( q=>pro_state_65, i=>nx652, ck=>
      conpro_system_clk);
   reg_pro_state_64 : sff1_x4 port map ( q=>pro_state_64, i=>nx642, ck=>
      conpro_system_clk);
   reg_pro_state_63 : sff1_x4 port map ( q=>pro_state_63, i=>nx632, ck=>
      conpro_system_clk);
   reg_pro_state_62 : sff1_x4 port map ( q=>pro_state_62, i=>nx622, ck=>
      conpro_system_clk);
   reg_pro_state_61 : sff1_x4 port map ( q=>pro_state_61, i=>nx612, ck=>
      conpro_system_clk);
   reg_pro_state_60 : sff1_x4 port map ( q=>pro_state_60, i=>nx602, ck=>
      conpro_system_clk);
   reg_pro_state_59 : sff1_x4 port map ( q=>pro_state_59, i=>nx592, ck=>
      conpro_system_clk);
   reg_pro_state_58 : sff1_x4 port map ( q=>pro_state_58, i=>nx582, ck=>
      conpro_system_clk);
   reg_pro_state_57 : sff1_x4 port map ( q=>pro_state_57, i=>nx572, ck=>
      conpro_system_clk);
   reg_pro_state_56 : sff1_x4 port map ( q=>pro_state_56, i=>nx562, ck=>
      conpro_system_clk);
   reg_pro_state_55 : sff1_x4 port map ( q=>pro_state_55, i=>nx552, ck=>
      conpro_system_clk);
   reg_pro_state_54 : sff1_x4 port map ( q=>pro_state_54, i=>nx542, ck=>
      conpro_system_clk);
   reg_pro_state_53 : sff1_x4 port map ( q=>pro_state_53, i=>nx532, ck=>
      conpro_system_clk);
   reg_pro_state_52 : sff1_x4 port map ( q=>pro_state_52, i=>nx522, ck=>
      conpro_system_clk);
   reg_pro_state_51 : sff1_x4 port map ( q=>pro_state_51, i=>nx512, ck=>
      conpro_system_clk);
   reg_pro_state_50 : sff1_x4 port map ( q=>pro_state_50, i=>nx502, ck=>
      conpro_system_clk);
   reg_pro_state_49 : sff1_x4 port map ( q=>pro_state_49, i=>nx492, ck=>
      conpro_system_clk);
   reg_pro_state_48 : sff1_x4 port map ( q=>pro_state_48, i=>nx482, ck=>
      conpro_system_clk);
   reg_pro_state_47 : sff1_x4 port map ( q=>pro_state_47, i=>nx472, ck=>
      conpro_system_clk);
   reg_pro_state_46 : sff1_x4 port map ( q=>pro_state_46, i=>nx462, ck=>
      conpro_system_clk);
   reg_pro_state_45 : sff1_x4 port map ( q=>pro_state_45, i=>nx452, ck=>
      conpro_system_clk);
   reg_pro_state_44 : sff1_x4 port map ( q=>pro_state_44, i=>nx442, ck=>
      conpro_system_clk);
   reg_pro_state_43 : sff1_x4 port map ( q=>pro_state_43, i=>nx432, ck=>
      conpro_system_clk);
   reg_pro_state_42 : sff1_x4 port map ( q=>pro_state_42, i=>nx422, ck=>
      conpro_system_clk);
   reg_pro_state_41 : sff1_x4 port map ( q=>pro_state_41, i=>nx412, ck=>
      conpro_system_clk);
   reg_pro_state_40 : sff1_x4 port map ( q=>pro_state_40, i=>nx402, ck=>
      conpro_system_clk);
   reg_pro_state_39 : sff1_x4 port map ( q=>pro_state_39, i=>nx392, ck=>
      conpro_system_clk);
   reg_pro_state_38 : sff1_x4 port map ( q=>pro_state_38, i=>nx382, ck=>
      conpro_system_clk);
   reg_pro_state_37 : sff1_x4 port map ( q=>pro_state_37, i=>nx372, ck=>
      conpro_system_clk);
   reg_pro_state_36 : sff1_x4 port map ( q=>pro_state_36, i=>nx362, ck=>
      conpro_system_clk);
   reg_pro_state_35 : sff1_x4 port map ( q=>pro_state_35, i=>nx352, ck=>
      conpro_system_clk);
   reg_pro_state_34 : sff1_x4 port map ( q=>pro_state_34, i=>nx342, ck=>
      conpro_system_clk);
   reg_pro_state_33 : sff1_x4 port map ( q=>pro_state_33, i=>nx332, ck=>
      conpro_system_clk);
   reg_pro_state_32 : sff1_x4 port map ( q=>pro_state_32, i=>nx322, ck=>
      conpro_system_clk);
   reg_pro_state_31 : sff1_x4 port map ( q=>pro_state_31, i=>nx312, ck=>
      conpro_system_clk);
   reg_pro_state_30 : sff1_x4 port map ( q=>pro_state_30, i=>nx302, ck=>
      conpro_system_clk);
   reg_pro_state_29 : sff1_x4 port map ( q=>pro_state_29, i=>nx292, ck=>
      conpro_system_clk);
   reg_pro_state_28 : sff1_x4 port map ( q=>pro_state_28, i=>nx282, ck=>
      conpro_system_clk);
   reg_pro_state_27 : sff1_x4 port map ( q=>pro_state_27, i=>nx272, ck=>
      conpro_system_clk);
   reg_pro_state_26 : sff1_x4 port map ( q=>pro_state_26, i=>nx262, ck=>
      conpro_system_clk);
   reg_pro_state_25 : sff1_x4 port map ( q=>pro_state_25, i=>nx252, ck=>
      conpro_system_clk);
   reg_pro_state_24 : sff1_x4 port map ( q=>pro_state_24, i=>nx242, ck=>
      conpro_system_clk);
   reg_pro_state_23 : sff1_x4 port map ( q=>pro_state_23, i=>nx232, ck=>
      conpro_system_clk);
   reg_pro_state_22 : sff1_x4 port map ( q=>pro_state_22, i=>nx222, ck=>
      conpro_system_clk);
   reg_pro_state_21 : sff1_x4 port map ( q=>pro_state_21, i=>nx212, ck=>
      conpro_system_clk);
   reg_pro_state_20 : sff1_x4 port map ( q=>pro_state_20, i=>nx202, ck=>
      conpro_system_clk);
   reg_pro_state_19 : sff1_x4 port map ( q=>pro_state_19, i=>nx192, ck=>
      conpro_system_clk);
   reg_pro_state_18 : sff1_x4 port map ( q=>pro_state_18, i=>nx182, ck=>
      conpro_system_clk);
   reg_pro_state_17 : sff1_x4 port map ( q=>pro_state_17, i=>nx172, ck=>
      conpro_system_clk);
   reg_pro_state_16 : sff1_x4 port map ( q=>pro_state_16, i=>nx162, ck=>
      conpro_system_clk);
   reg_pro_state_15 : sff1_x4 port map ( q=>pro_state_15, i=>nx152, ck=>
      conpro_system_clk);
   reg_pro_state_14 : sff1_x4 port map ( q=>pro_state_14, i=>nx142, ck=>
      conpro_system_clk);
   reg_pro_state_13 : sff1_x4 port map ( q=>pro_state_13, i=>nx132, ck=>
      conpro_system_clk);
   reg_pro_state_12 : sff1_x4 port map ( q=>pro_state_12, i=>nx122, ck=>
      conpro_system_clk);
   reg_pro_state_11 : sff1_x4 port map ( q=>pro_state_11, i=>nx112, ck=>
      conpro_system_clk);
   reg_pro_state_10 : sff1_x4 port map ( q=>pro_state_10, i=>nx102, ck=>
      conpro_system_clk);
   reg_pro_state_9 : sff1_x4 port map ( q=>pro_state_9, i=>nx92, ck=>
      conpro_system_clk);
   reg_pro_state_8 : sff1_x4 port map ( q=>pro_state_8, i=>nx82, ck=>
      conpro_system_clk);
   reg_pro_state_7 : sff1_x4 port map ( q=>pro_state_7, i=>nx72, ck=>
      conpro_system_clk);
   reg_pro_state_6 : sff1_x4 port map ( q=>pro_state_6, i=>nx62, ck=>
      conpro_system_clk);
   reg_pro_state_5 : sff1_x4 port map ( q=>pro_state_5, i=>nx52, ck=>
      conpro_system_clk);
   reg_pro_state_4 : sff1_x4 port map ( q=>pro_state_4, i=>nx42, ck=>
      conpro_system_clk);
   reg_pro_state_3 : sff1_x4 port map ( q=>pro_state_3, i=>nx32, ck=>
      conpro_system_clk);
   ix33 : an12_x1 port map ( q=>nx32, i0=>nx3589, i1=>pro_state_2);
   reg_pro_state_2 : sff1_x4 port map ( q=>pro_state_2, i=>nx22, ck=>
      conpro_system_clk);
   reg_pro_state_1 : sff1_x4 port map ( q=>pro_state_1, i=>nx12, ck=>
      conpro_system_clk);
   reg_pro_state_0 : sff1_x4 port map ( q=>pro_state_0, i=>nx3589, ck=>
      conpro_system_clk);
   reg_pl : sff2_x4 port map ( q=>pl, i0=>nx3611, i1=>nx1734, cmd=>nx706, ck
      =>conpro_system_clk);
   ix1735 : no2_x1 port map ( nq=>nx1734, i0=>conpro_system_reset, i1=>
      nx3346);
   ix3347 : no4_x1 port map ( nq=>nx3346, i0=>nx1726, i1=>nx1472, i2=>nx1216, 
      i3=>nx962);
   ix1727 : na4_x1 port map ( nq=>nx1726, i0=>nx3349, i1=>nx3364, i2=>nx3378, 
      i3=>nx3392);
   ix3350 : noa2a2a2a24_x1 port map ( nq=>nx3349, i0=>pro_state_66, i1=>
      nx1716, i2=>pro_state_65, i3=>nx1702, i4=>pro_state_64, i5=>nx1686, i6
      =>pro_state_63, i7=>nx1672);
   ix1717 : xr2_x1 port map ( q=>nx1716, i0=>nx3611, i1=>xl_63);
   reg_xl_63 : sff2_x4 port map ( q=>xl_63, i0=>xl_63, i1=>nx1708, cmd=>
      nx3619, ck=>conpro_system_clk);
   ix1709 : an12_x1 port map ( q=>nx1708, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(63));
   ix1703 : xr2_x1 port map ( q=>nx1702, i0=>nx3611, i1=>xl_62);
   reg_xl_62 : sff2_x4 port map ( q=>xl_62, i0=>xl_62, i1=>nx1694, cmd=>
      nx3619, ck=>conpro_system_clk);
   ix1695 : an12_x1 port map ( q=>nx1694, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(62));
   ix1687 : xr2_x1 port map ( q=>nx1686, i0=>nx3611, i1=>xl_61);
   reg_xl_61 : sff2_x4 port map ( q=>xl_61, i0=>xl_61, i1=>nx1678, cmd=>
      nx3619, ck=>conpro_system_clk);
   ix1679 : an12_x1 port map ( q=>nx1678, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(61));
   ix1673 : xr2_x1 port map ( q=>nx1672, i0=>nx3611, i1=>xl_60);
   reg_xl_60 : sff2_x4 port map ( q=>xl_60, i0=>xl_60, i1=>nx1664, cmd=>
      nx3619, ck=>conpro_system_clk);
   ix1665 : an12_x1 port map ( q=>nx1664, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(60));
   ix3365 : noa2a2a2a24_x1 port map ( nq=>nx3364, i0=>pro_state_62, i1=>
      nx1654, i2=>pro_state_61, i3=>nx1640, i4=>pro_state_60, i5=>nx1624, i6
      =>pro_state_59, i7=>nx1610);
   ix1655 : xr2_x1 port map ( q=>nx1654, i0=>nx3611, i1=>xl_59);
   reg_xl_59 : sff2_x4 port map ( q=>xl_59, i0=>xl_59, i1=>nx1646, cmd=>
      nx3621, ck=>conpro_system_clk);
   ix1647 : an12_x1 port map ( q=>nx1646, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(59));
   ix1641 : xr2_x1 port map ( q=>nx1640, i0=>nx3611, i1=>xl_58);
   reg_xl_58 : sff2_x4 port map ( q=>xl_58, i0=>xl_58, i1=>nx1632, cmd=>
      nx3621, ck=>conpro_system_clk);
   ix1633 : an12_x1 port map ( q=>nx1632, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(58));
   ix1625 : xr2_x1 port map ( q=>nx1624, i0=>nx3611, i1=>xl_57);
   reg_xl_57 : sff2_x4 port map ( q=>xl_57, i0=>xl_57, i1=>nx1616, cmd=>
      nx3621, ck=>conpro_system_clk);
   ix1617 : an12_x1 port map ( q=>nx1616, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(57));
   ix1611 : xr2_x1 port map ( q=>nx1610, i0=>nx3611, i1=>xl_56);
   reg_xl_56 : sff2_x4 port map ( q=>xl_56, i0=>xl_56, i1=>nx1602, cmd=>
      nx3621, ck=>conpro_system_clk);
   ix1603 : an12_x1 port map ( q=>nx1602, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(56));
   ix3379 : noa2a2a2a24_x1 port map ( nq=>nx3378, i0=>pro_state_58, i1=>
      nx1590, i2=>pro_state_57, i3=>nx1576, i4=>pro_state_56, i5=>nx1560, i6
      =>pro_state_55, i7=>nx1546);
   ix1591 : xr2_x1 port map ( q=>nx1590, i0=>nx3611, i1=>xl_55);
   reg_xl_55 : sff2_x4 port map ( q=>xl_55, i0=>xl_55, i1=>nx1582, cmd=>
      nx3623, ck=>conpro_system_clk);
   ix1583 : an12_x1 port map ( q=>nx1582, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(55));
   ix1577 : xr2_x1 port map ( q=>nx1576, i0=>nx3611, i1=>xl_54);
   reg_xl_54 : sff2_x4 port map ( q=>xl_54, i0=>xl_54, i1=>nx1568, cmd=>
      nx3623, ck=>conpro_system_clk);
   ix1569 : an12_x1 port map ( q=>nx1568, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(54));
   ix1561 : xr2_x1 port map ( q=>nx1560, i0=>nx3611, i1=>xl_53);
   reg_xl_53 : sff2_x4 port map ( q=>xl_53, i0=>xl_53, i1=>nx1552, cmd=>
      nx3623, ck=>conpro_system_clk);
   ix1553 : an12_x1 port map ( q=>nx1552, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(53));
   ix1547 : xr2_x1 port map ( q=>nx1546, i0=>nx3611, i1=>xl_52);
   reg_xl_52 : sff2_x4 port map ( q=>xl_52, i0=>xl_52, i1=>nx1538, cmd=>
      nx3623, ck=>conpro_system_clk);
   ix1539 : an12_x1 port map ( q=>nx1538, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(52));
   ix3393 : noa2a2a2a24_x1 port map ( nq=>nx3392, i0=>pro_state_54, i1=>
      nx1528, i2=>pro_state_53, i3=>nx1514, i4=>pro_state_52, i5=>nx1498, i6
      =>pro_state_51, i7=>nx1484);
   ix1529 : xr2_x1 port map ( q=>nx1528, i0=>nx3611, i1=>xl_51);
   reg_xl_51 : sff2_x4 port map ( q=>xl_51, i0=>xl_51, i1=>nx1520, cmd=>
      nx3625, ck=>conpro_system_clk);
   ix1521 : an12_x1 port map ( q=>nx1520, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(51));
   ix1515 : xr2_x1 port map ( q=>nx1514, i0=>nx3611, i1=>xl_50);
   reg_xl_50 : sff2_x4 port map ( q=>xl_50, i0=>xl_50, i1=>nx1506, cmd=>
      nx3625, ck=>conpro_system_clk);
   ix1507 : an12_x1 port map ( q=>nx1506, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(50));
   ix1499 : xr2_x1 port map ( q=>nx1498, i0=>nx3613, i1=>xl_49);
   reg_xl_49 : sff2_x4 port map ( q=>xl_49, i0=>xl_49, i1=>nx1490, cmd=>
      nx3625, ck=>conpro_system_clk);
   ix1491 : an12_x1 port map ( q=>nx1490, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(49));
   ix1485 : xr2_x1 port map ( q=>nx1484, i0=>nx3613, i1=>xl_48);
   reg_xl_48 : sff2_x4 port map ( q=>xl_48, i0=>xl_48, i1=>nx1476, cmd=>
      nx3625, ck=>conpro_system_clk);
   ix1477 : an12_x1 port map ( q=>nx1476, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(48));
   ix1473 : na4_x1 port map ( nq=>nx1472, i0=>nx3407, i1=>nx3421, i2=>nx3435, 
      i3=>nx3449);
   ix3408 : noa2a2a2a24_x1 port map ( nq=>nx3407, i0=>pro_state_50, i1=>
      nx1462, i2=>pro_state_49, i3=>nx1448, i4=>pro_state_48, i5=>nx1432, i6
      =>pro_state_47, i7=>nx1418);
   ix1463 : xr2_x1 port map ( q=>nx1462, i0=>nx3613, i1=>xl_47);
   reg_xl_47 : sff2_x4 port map ( q=>xl_47, i0=>xl_47, i1=>nx1454, cmd=>
      nx3627, ck=>conpro_system_clk);
   ix1455 : an12_x1 port map ( q=>nx1454, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(47));
   ix1449 : xr2_x1 port map ( q=>nx1448, i0=>nx3613, i1=>xl_46);
   reg_xl_46 : sff2_x4 port map ( q=>xl_46, i0=>xl_46, i1=>nx1440, cmd=>
      nx3627, ck=>conpro_system_clk);
   ix1441 : an12_x1 port map ( q=>nx1440, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(46));
   ix1433 : xr2_x1 port map ( q=>nx1432, i0=>nx3613, i1=>xl_45);
   reg_xl_45 : sff2_x4 port map ( q=>xl_45, i0=>xl_45, i1=>nx1424, cmd=>
      nx3627, ck=>conpro_system_clk);
   ix1425 : an12_x1 port map ( q=>nx1424, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(45));
   ix1419 : xr2_x1 port map ( q=>nx1418, i0=>nx3613, i1=>xl_44);
   reg_xl_44 : sff2_x4 port map ( q=>xl_44, i0=>xl_44, i1=>nx1410, cmd=>
      nx3627, ck=>conpro_system_clk);
   ix1411 : an12_x1 port map ( q=>nx1410, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(44));
   ix3422 : noa2a2a2a24_x1 port map ( nq=>nx3421, i0=>pro_state_46, i1=>
      nx1400, i2=>pro_state_45, i3=>nx1386, i4=>pro_state_44, i5=>nx1370, i6
      =>pro_state_43, i7=>nx1356);
   ix1401 : xr2_x1 port map ( q=>nx1400, i0=>nx3613, i1=>xl_43);
   reg_xl_43 : sff2_x4 port map ( q=>xl_43, i0=>xl_43, i1=>nx1392, cmd=>
      nx3629, ck=>conpro_system_clk);
   ix1393 : an12_x1 port map ( q=>nx1392, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(43));
   ix1387 : xr2_x1 port map ( q=>nx1386, i0=>nx3613, i1=>xl_42);
   reg_xl_42 : sff2_x4 port map ( q=>xl_42, i0=>xl_42, i1=>nx1378, cmd=>
      nx3629, ck=>conpro_system_clk);
   ix1379 : an12_x1 port map ( q=>nx1378, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(42));
   ix1371 : xr2_x1 port map ( q=>nx1370, i0=>nx3613, i1=>xl_41);
   reg_xl_41 : sff2_x4 port map ( q=>xl_41, i0=>xl_41, i1=>nx1362, cmd=>
      nx3629, ck=>conpro_system_clk);
   ix1363 : an12_x1 port map ( q=>nx1362, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(41));
   ix1357 : xr2_x1 port map ( q=>nx1356, i0=>nx3613, i1=>xl_40);
   reg_xl_40 : sff2_x4 port map ( q=>xl_40, i0=>xl_40, i1=>nx1348, cmd=>
      nx3629, ck=>conpro_system_clk);
   ix1349 : an12_x1 port map ( q=>nx1348, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(40));
   ix3436 : noa2a2a2a24_x1 port map ( nq=>nx3435, i0=>pro_state_42, i1=>
      nx1336, i2=>pro_state_41, i3=>nx1322, i4=>pro_state_40, i5=>nx1306, i6
      =>pro_state_39, i7=>nx1292);
   ix1337 : xr2_x1 port map ( q=>nx1336, i0=>nx3613, i1=>xl_39);
   reg_xl_39 : sff2_x4 port map ( q=>xl_39, i0=>xl_39, i1=>nx1328, cmd=>
      nx3631, ck=>conpro_system_clk);
   ix1329 : an12_x1 port map ( q=>nx1328, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(39));
   ix1323 : xr2_x1 port map ( q=>nx1322, i0=>nx3613, i1=>xl_38);
   reg_xl_38 : sff2_x4 port map ( q=>xl_38, i0=>xl_38, i1=>nx1314, cmd=>
      nx3631, ck=>conpro_system_clk);
   ix1315 : an12_x1 port map ( q=>nx1314, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(38));
   ix1307 : xr2_x1 port map ( q=>nx1306, i0=>nx3613, i1=>xl_37);
   reg_xl_37 : sff2_x4 port map ( q=>xl_37, i0=>xl_37, i1=>nx1298, cmd=>
      nx3631, ck=>conpro_system_clk);
   ix1299 : an12_x1 port map ( q=>nx1298, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(37));
   ix1293 : xr2_x1 port map ( q=>nx1292, i0=>nx3613, i1=>xl_36);
   reg_xl_36 : sff2_x4 port map ( q=>xl_36, i0=>xl_36, i1=>nx1284, cmd=>
      nx3631, ck=>conpro_system_clk);
   ix1285 : an12_x1 port map ( q=>nx1284, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(36));
   ix3450 : noa2a2a2a24_x1 port map ( nq=>nx3449, i0=>pro_state_38, i1=>
      nx1274, i2=>pro_state_37, i3=>nx1260, i4=>pro_state_36, i5=>nx1244, i6
      =>pro_state_35, i7=>nx1230);
   ix1275 : xr2_x1 port map ( q=>nx1274, i0=>nx3615, i1=>xl_35);
   reg_xl_35 : sff2_x4 port map ( q=>xl_35, i0=>xl_35, i1=>nx1266, cmd=>
      nx3633, ck=>conpro_system_clk);
   ix1267 : an12_x1 port map ( q=>nx1266, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(35));
   ix1261 : xr2_x1 port map ( q=>nx1260, i0=>nx3615, i1=>xl_34);
   reg_xl_34 : sff2_x4 port map ( q=>xl_34, i0=>xl_34, i1=>nx1252, cmd=>
      nx3633, ck=>conpro_system_clk);
   ix1253 : an12_x1 port map ( q=>nx1252, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(34));
   ix1245 : xr2_x1 port map ( q=>nx1244, i0=>nx3615, i1=>xl_33);
   reg_xl_33 : sff2_x4 port map ( q=>xl_33, i0=>xl_33, i1=>nx1236, cmd=>
      nx3633, ck=>conpro_system_clk);
   ix1237 : an12_x1 port map ( q=>nx1236, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(33));
   ix1231 : xr2_x1 port map ( q=>nx1230, i0=>nx3615, i1=>xl_32);
   reg_xl_32 : sff2_x4 port map ( q=>xl_32, i0=>xl_32, i1=>nx1222, cmd=>
      nx3633, ck=>conpro_system_clk);
   ix1223 : an12_x1 port map ( q=>nx1222, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(32));
   ix1217 : na4_x1 port map ( nq=>nx1216, i0=>nx3464, i1=>nx3478, i2=>nx3492, 
      i3=>nx3506);
   ix3465 : noa2a2a2a24_x1 port map ( nq=>nx3464, i0=>pro_state_34, i1=>
      nx1206, i2=>pro_state_33, i3=>nx1192, i4=>pro_state_32, i5=>nx1176, i6
      =>pro_state_31, i7=>nx1162);
   ix1207 : xr2_x1 port map ( q=>nx1206, i0=>nx3615, i1=>xl_31);
   reg_xl_31 : sff2_x4 port map ( q=>xl_31, i0=>xl_31, i1=>nx1198, cmd=>
      nx3635, ck=>conpro_system_clk);
   ix1199 : an12_x1 port map ( q=>nx1198, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(31));
   ix1193 : xr2_x1 port map ( q=>nx1192, i0=>nx3615, i1=>xl_30);
   reg_xl_30 : sff2_x4 port map ( q=>xl_30, i0=>xl_30, i1=>nx1184, cmd=>
      nx3635, ck=>conpro_system_clk);
   ix1185 : an12_x1 port map ( q=>nx1184, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(30));
   ix1177 : xr2_x1 port map ( q=>nx1176, i0=>nx3615, i1=>xl_29);
   reg_xl_29 : sff2_x4 port map ( q=>xl_29, i0=>xl_29, i1=>nx1168, cmd=>
      nx3635, ck=>conpro_system_clk);
   ix1169 : an12_x1 port map ( q=>nx1168, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(29));
   ix1163 : xr2_x1 port map ( q=>nx1162, i0=>nx3615, i1=>xl_28);
   reg_xl_28 : sff2_x4 port map ( q=>xl_28, i0=>xl_28, i1=>nx1154, cmd=>
      nx3635, ck=>conpro_system_clk);
   ix1155 : an12_x1 port map ( q=>nx1154, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(28));
   ix3479 : noa2a2a2a24_x1 port map ( nq=>nx3478, i0=>pro_state_30, i1=>
      nx1144, i2=>pro_state_29, i3=>nx1130, i4=>pro_state_28, i5=>nx1114, i6
      =>pro_state_27, i7=>nx1100);
   ix1145 : xr2_x1 port map ( q=>nx1144, i0=>nx3615, i1=>xl_27);
   reg_xl_27 : sff2_x4 port map ( q=>xl_27, i0=>xl_27, i1=>nx1136, cmd=>
      nx3637, ck=>conpro_system_clk);
   ix1137 : an12_x1 port map ( q=>nx1136, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(27));
   ix1131 : xr2_x1 port map ( q=>nx1130, i0=>nx3615, i1=>xl_26);
   reg_xl_26 : sff2_x4 port map ( q=>xl_26, i0=>xl_26, i1=>nx1122, cmd=>
      nx3637, ck=>conpro_system_clk);
   ix1123 : an12_x1 port map ( q=>nx1122, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(26));
   ix1115 : xr2_x1 port map ( q=>nx1114, i0=>nx3615, i1=>xl_25);
   reg_xl_25 : sff2_x4 port map ( q=>xl_25, i0=>xl_25, i1=>nx1106, cmd=>
      nx3637, ck=>conpro_system_clk);
   ix1107 : an12_x1 port map ( q=>nx1106, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(25));
   ix1101 : xr2_x1 port map ( q=>nx1100, i0=>nx3615, i1=>xl_24);
   reg_xl_24 : sff2_x4 port map ( q=>xl_24, i0=>xl_24, i1=>nx1092, cmd=>
      nx3637, ck=>conpro_system_clk);
   ix1093 : an12_x1 port map ( q=>nx1092, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(24));
   ix3493 : noa2a2a2a24_x1 port map ( nq=>nx3492, i0=>pro_state_26, i1=>
      nx1080, i2=>pro_state_25, i3=>nx1066, i4=>pro_state_24, i5=>nx1050, i6
      =>pro_state_23, i7=>nx1036);
   ix1081 : xr2_x1 port map ( q=>nx1080, i0=>nx3615, i1=>xl_23);
   reg_xl_23 : sff2_x4 port map ( q=>xl_23, i0=>xl_23, i1=>nx1072, cmd=>
      nx3639, ck=>conpro_system_clk);
   ix1073 : an12_x1 port map ( q=>nx1072, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(23));
   ix1067 : xr2_x1 port map ( q=>nx1066, i0=>nx3615, i1=>xl_22);
   reg_xl_22 : sff2_x4 port map ( q=>xl_22, i0=>xl_22, i1=>nx1058, cmd=>
      nx3639, ck=>conpro_system_clk);
   ix1059 : an12_x1 port map ( q=>nx1058, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(22));
   ix1051 : xr2_x1 port map ( q=>nx1050, i0=>nx3617, i1=>xl_21);
   reg_xl_21 : sff2_x4 port map ( q=>xl_21, i0=>xl_21, i1=>nx1042, cmd=>
      nx3639, ck=>conpro_system_clk);
   ix1043 : an12_x1 port map ( q=>nx1042, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(21));
   ix1037 : xr2_x1 port map ( q=>nx1036, i0=>nx3617, i1=>xl_20);
   reg_xl_20 : sff2_x4 port map ( q=>xl_20, i0=>xl_20, i1=>nx1028, cmd=>
      nx3639, ck=>conpro_system_clk);
   ix1029 : an12_x1 port map ( q=>nx1028, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(20));
   ix3507 : noa2a2a2a24_x1 port map ( nq=>nx3506, i0=>pro_state_22, i1=>
      nx1018, i2=>pro_state_21, i3=>nx1004, i4=>pro_state_20, i5=>nx988, i6
      =>pro_state_19, i7=>nx974);
   ix1019 : xr2_x1 port map ( q=>nx1018, i0=>nx3617, i1=>xl_19);
   reg_xl_19 : sff2_x4 port map ( q=>xl_19, i0=>xl_19, i1=>nx1010, cmd=>
      nx3641, ck=>conpro_system_clk);
   ix1011 : an12_x1 port map ( q=>nx1010, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(19));
   ix1005 : xr2_x1 port map ( q=>nx1004, i0=>nx3617, i1=>xl_18);
   reg_xl_18 : sff2_x4 port map ( q=>xl_18, i0=>xl_18, i1=>nx996, cmd=>
      nx3641, ck=>conpro_system_clk);
   ix997 : an12_x1 port map ( q=>nx996, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(18));
   ix989 : xr2_x1 port map ( q=>nx988, i0=>nx3617, i1=>xl_17);
   reg_xl_17 : sff2_x4 port map ( q=>xl_17, i0=>xl_17, i1=>nx980, cmd=>
      nx3641, ck=>conpro_system_clk);
   ix981 : an12_x1 port map ( q=>nx980, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(17));
   ix975 : xr2_x1 port map ( q=>nx974, i0=>nx3617, i1=>xl_16);
   reg_xl_16 : sff2_x4 port map ( q=>xl_16, i0=>xl_16, i1=>nx966, cmd=>
      nx3641, ck=>conpro_system_clk);
   ix967 : an12_x1 port map ( q=>nx966, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(16));
   ix963 : na4_x1 port map ( nq=>nx962, i0=>nx3521, i1=>nx3535, i2=>nx3549, 
      i3=>nx3563);
   ix3522 : noa2a2a2a24_x1 port map ( nq=>nx3521, i0=>pro_state_18, i1=>
      nx952, i2=>pro_state_17, i3=>nx938, i4=>pro_state_16, i5=>nx922, i6=>
      pro_state_15, i7=>nx908);
   ix953 : xr2_x1 port map ( q=>nx952, i0=>nx3617, i1=>xl_15);
   reg_xl_15 : sff2_x4 port map ( q=>xl_15, i0=>xl_15, i1=>nx944, cmd=>
      nx3643, ck=>conpro_system_clk);
   ix945 : an12_x1 port map ( q=>nx944, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(15));
   ix939 : xr2_x1 port map ( q=>nx938, i0=>nx3617, i1=>xl_14);
   reg_xl_14 : sff2_x4 port map ( q=>xl_14, i0=>xl_14, i1=>nx930, cmd=>
      nx3643, ck=>conpro_system_clk);
   ix931 : an12_x1 port map ( q=>nx930, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(14));
   ix923 : xr2_x1 port map ( q=>nx922, i0=>nx3617, i1=>xl_13);
   reg_xl_13 : sff2_x4 port map ( q=>xl_13, i0=>xl_13, i1=>nx914, cmd=>
      nx3643, ck=>conpro_system_clk);
   ix915 : an12_x1 port map ( q=>nx914, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(13));
   ix909 : xr2_x1 port map ( q=>nx908, i0=>nx3617, i1=>xl_12);
   reg_xl_12 : sff2_x4 port map ( q=>xl_12, i0=>xl_12, i1=>nx900, cmd=>
      nx3643, ck=>conpro_system_clk);
   ix901 : an12_x1 port map ( q=>nx900, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(12));
   ix3536 : noa2a2a2a24_x1 port map ( nq=>nx3535, i0=>pro_state_14, i1=>
      nx890, i2=>pro_state_13, i3=>nx876, i4=>pro_state_12, i5=>nx860, i6=>
      pro_state_11, i7=>nx846);
   ix891 : xr2_x1 port map ( q=>nx890, i0=>nx3617, i1=>xl_11);
   reg_xl_11 : sff2_x4 port map ( q=>xl_11, i0=>xl_11, i1=>nx882, cmd=>
      nx3645, ck=>conpro_system_clk);
   ix883 : an12_x1 port map ( q=>nx882, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(11));
   ix877 : xr2_x1 port map ( q=>nx876, i0=>nx3617, i1=>xl_10);
   reg_xl_10 : sff2_x4 port map ( q=>xl_10, i0=>xl_10, i1=>nx868, cmd=>
      nx3645, ck=>conpro_system_clk);
   ix869 : an12_x1 port map ( q=>nx868, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(10));
   ix861 : xr2_x1 port map ( q=>nx860, i0=>nx3617, i1=>xl_9);
   reg_xl_9 : sff2_x4 port map ( q=>xl_9, i0=>xl_9, i1=>nx852, cmd=>nx3645, 
      ck=>conpro_system_clk);
   ix853 : an12_x1 port map ( q=>nx852, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(9));
   ix847 : xr2_x1 port map ( q=>nx846, i0=>nx3617, i1=>xl_8);
   reg_xl_8 : sff2_x4 port map ( q=>xl_8, i0=>xl_8, i1=>nx838, cmd=>nx3645, 
      ck=>conpro_system_clk);
   ix839 : an12_x1 port map ( q=>nx838, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(8));
   ix3550 : noa2a2a2a24_x1 port map ( nq=>nx3549, i0=>pro_state_10, i1=>
      nx826, i2=>pro_state_9, i3=>nx812, i4=>pro_state_8, i5=>nx796, i6=>
      pro_state_7, i7=>nx782);
   ix827 : xr2_x1 port map ( q=>nx826, i0=>pl, i1=>xl_7);
   reg_xl_7 : sff2_x4 port map ( q=>xl_7, i0=>xl_7, i1=>nx818, cmd=>nx3647, 
      ck=>conpro_system_clk);
   ix819 : an12_x1 port map ( q=>nx818, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(7));
   ix813 : xr2_x1 port map ( q=>nx812, i0=>pl, i1=>xl_6);
   reg_xl_6 : sff2_x4 port map ( q=>xl_6, i0=>xl_6, i1=>nx804, cmd=>nx3647, 
      ck=>conpro_system_clk);
   ix805 : an12_x1 port map ( q=>nx804, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(6));
   ix797 : xr2_x1 port map ( q=>nx796, i0=>pl, i1=>xl_5);
   reg_xl_5 : sff2_x4 port map ( q=>xl_5, i0=>xl_5, i1=>nx788, cmd=>nx3647, 
      ck=>conpro_system_clk);
   ix789 : an12_x1 port map ( q=>nx788, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(5));
   ix783 : xr2_x1 port map ( q=>nx782, i0=>pl, i1=>xl_4);
   reg_xl_4 : sff2_x4 port map ( q=>xl_4, i0=>xl_4, i1=>nx774, cmd=>nx3647, 
      ck=>conpro_system_clk);
   ix775 : an12_x1 port map ( q=>nx774, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(4));
   ix3564 : noa2a2a2a24_x1 port map ( nq=>nx3563, i0=>pro_state_6, i1=>nx764, 
      i2=>pro_state_5, i3=>nx750, i4=>pro_state_4, i5=>nx734, i6=>
      pro_state_3, i7=>nx720);
   ix765 : xr2_x1 port map ( q=>nx764, i0=>pl, i1=>xl_3);
   reg_xl_3 : sff2_x4 port map ( q=>xl_3, i0=>xl_3, i1=>nx756, cmd=>nx708, 
      ck=>conpro_system_clk);
   ix757 : an12_x1 port map ( q=>nx756, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(3));
   ix751 : xr2_x1 port map ( q=>nx750, i0=>pl, i1=>xl_2);
   reg_xl_2 : sff2_x4 port map ( q=>xl_2, i0=>xl_2, i1=>nx742, cmd=>nx708, 
      ck=>conpro_system_clk);
   ix743 : an12_x1 port map ( q=>nx742, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(2));
   ix735 : xr2_x1 port map ( q=>nx734, i0=>pl, i1=>xl_1);
   reg_xl_1 : sff2_x4 port map ( q=>xl_1, i0=>xl_1, i1=>nx726, cmd=>nx708, 
      ck=>conpro_system_clk);
   ix727 : an12_x1 port map ( q=>nx726, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(1));
   ix721 : xr2_x1 port map ( q=>nx720, i0=>pl, i1=>xl_0);
   reg_xl_0 : sff2_x4 port map ( q=>xl_0, i0=>xl_0, i1=>nx712, cmd=>nx708, 
      ck=>conpro_system_clk);
   ix713 : an12_x1 port map ( q=>nx712, i0=>conpro_system_reset, i1=>
      REG_ARG_FUN_parity3_x_RD(0));
   ix3579 : o4_x2 port map ( q=>nx3578, i0=>PRO_FUN_parity3_END_EXMPLR, i1=>
      REG_RET_FUN_parity3_p_WE_EXMPLR, i2=>pro_state_1, i3=>pro_state_0);
   reg_pro_state_68 : sff1_x4 port map ( q=>PRO_FUN_parity3_END_EXMPLR, i=>
      nx684, ck=>conpro_system_clk);
   ix685 : ao22_x2 port map ( q=>nx684, i0=>REG_RET_FUN_parity3_p_WE_EXMPLR, 
      i1=>PRO_FUN_parity3_END_EXMPLR, i2=>nx3582);
   ix3583 : inv_x1 port map ( nq=>nx3582, i=>nx2);
   reg_pl_rep_1 : sff2_x4 port map ( q=>nx3611, i0=>pl, i1=>nx1734, cmd=>
      nx706, ck=>conpro_system_clk);
   reg_pl_rep_2 : sff2_x4 port map ( q=>nx3613, i0=>nx3611, i1=>nx1734, cmd
      =>nx706, ck=>conpro_system_clk);
   reg_pl_rep_3 : sff2_x4 port map ( q=>nx3615, i0=>nx3611, i1=>nx1734, cmd
      =>nx706, ck=>conpro_system_clk);
   reg_pl_rep_4 : sff2_x4 port map ( q=>nx3617, i0=>nx3611, i1=>nx1734, cmd
      =>nx706, ck=>conpro_system_clk);
   ix673 : an12_x1 port map ( q=>nx672, i0=>nx2, i1=>pro_state_66);
   ix663 : an12_x1 port map ( q=>nx662, i0=>nx2, i1=>pro_state_65);
   ix653 : an12_x1 port map ( q=>nx652, i0=>nx3609, i1=>pro_state_64);
   ix643 : an12_x1 port map ( q=>nx642, i0=>nx3609, i1=>pro_state_63);
   ix633 : an12_x1 port map ( q=>nx632, i0=>nx3609, i1=>pro_state_62);
   ix623 : an12_x1 port map ( q=>nx622, i0=>nx3609, i1=>pro_state_61);
   ix613 : an12_x1 port map ( q=>nx612, i0=>nx3609, i1=>pro_state_60);
   ix603 : an12_x1 port map ( q=>nx602, i0=>nx3609, i1=>pro_state_59);
   ix593 : an12_x1 port map ( q=>nx592, i0=>nx3607, i1=>pro_state_58);
   ix583 : an12_x1 port map ( q=>nx582, i0=>nx3607, i1=>pro_state_57);
   ix573 : an12_x1 port map ( q=>nx572, i0=>nx3607, i1=>pro_state_56);
   ix563 : an12_x1 port map ( q=>nx562, i0=>nx3607, i1=>pro_state_55);
   ix553 : an12_x1 port map ( q=>nx552, i0=>nx3607, i1=>pro_state_54);
   ix543 : an12_x1 port map ( q=>nx542, i0=>nx3607, i1=>pro_state_53);
   ix533 : an12_x1 port map ( q=>nx532, i0=>nx3605, i1=>pro_state_52);
   ix523 : an12_x1 port map ( q=>nx522, i0=>nx3605, i1=>pro_state_51);
   ix513 : an12_x1 port map ( q=>nx512, i0=>nx3605, i1=>pro_state_50);
   ix503 : an12_x1 port map ( q=>nx502, i0=>nx3605, i1=>pro_state_49);
   ix493 : an12_x1 port map ( q=>nx492, i0=>nx3605, i1=>pro_state_48);
   ix483 : an12_x1 port map ( q=>nx482, i0=>nx3605, i1=>pro_state_47);
   ix473 : an12_x1 port map ( q=>nx472, i0=>nx3603, i1=>pro_state_46);
   ix463 : an12_x1 port map ( q=>nx462, i0=>nx3603, i1=>pro_state_45);
   ix453 : an12_x1 port map ( q=>nx452, i0=>nx3603, i1=>pro_state_44);
   ix443 : an12_x1 port map ( q=>nx442, i0=>nx3603, i1=>pro_state_43);
   ix433 : an12_x1 port map ( q=>nx432, i0=>nx3603, i1=>pro_state_42);
   ix423 : an12_x1 port map ( q=>nx422, i0=>nx3603, i1=>pro_state_41);
   ix413 : an12_x1 port map ( q=>nx412, i0=>nx3601, i1=>pro_state_40);
   ix403 : an12_x1 port map ( q=>nx402, i0=>nx3601, i1=>pro_state_39);
   ix393 : an12_x1 port map ( q=>nx392, i0=>nx3601, i1=>pro_state_38);
   ix383 : an12_x1 port map ( q=>nx382, i0=>nx3601, i1=>pro_state_37);
   ix373 : an12_x1 port map ( q=>nx372, i0=>nx3601, i1=>pro_state_36);
   ix363 : an12_x1 port map ( q=>nx362, i0=>nx3601, i1=>pro_state_35);
   ix353 : an12_x1 port map ( q=>nx352, i0=>nx3599, i1=>pro_state_34);
   ix343 : an12_x1 port map ( q=>nx342, i0=>nx3599, i1=>pro_state_33);
   ix333 : an12_x1 port map ( q=>nx332, i0=>nx3599, i1=>pro_state_32);
   ix323 : an12_x1 port map ( q=>nx322, i0=>nx3599, i1=>pro_state_31);
   ix313 : an12_x1 port map ( q=>nx312, i0=>nx3599, i1=>pro_state_30);
   ix303 : an12_x1 port map ( q=>nx302, i0=>nx3599, i1=>pro_state_29);
   ix293 : an12_x1 port map ( q=>nx292, i0=>nx3597, i1=>pro_state_28);
   ix283 : an12_x1 port map ( q=>nx282, i0=>nx3597, i1=>pro_state_27);
   ix273 : an12_x1 port map ( q=>nx272, i0=>nx3597, i1=>pro_state_26);
   ix263 : an12_x1 port map ( q=>nx262, i0=>nx3597, i1=>pro_state_25);
   ix253 : an12_x1 port map ( q=>nx252, i0=>nx3597, i1=>pro_state_24);
   ix243 : an12_x1 port map ( q=>nx242, i0=>nx3597, i1=>pro_state_23);
   ix233 : an12_x1 port map ( q=>nx232, i0=>nx3595, i1=>pro_state_22);
   ix223 : an12_x1 port map ( q=>nx222, i0=>nx3595, i1=>pro_state_21);
   ix213 : an12_x1 port map ( q=>nx212, i0=>nx3595, i1=>pro_state_20);
   ix203 : an12_x1 port map ( q=>nx202, i0=>nx3595, i1=>pro_state_19);
   ix193 : an12_x1 port map ( q=>nx192, i0=>nx3595, i1=>pro_state_18);
   ix183 : an12_x1 port map ( q=>nx182, i0=>nx3595, i1=>pro_state_17);
   ix173 : an12_x1 port map ( q=>nx172, i0=>nx3593, i1=>pro_state_16);
   ix163 : an12_x1 port map ( q=>nx162, i0=>nx3593, i1=>pro_state_15);
   ix153 : an12_x1 port map ( q=>nx152, i0=>nx3593, i1=>pro_state_14);
   ix143 : an12_x1 port map ( q=>nx142, i0=>nx3593, i1=>pro_state_13);
   ix133 : an12_x1 port map ( q=>nx132, i0=>nx3593, i1=>pro_state_12);
   ix123 : an12_x1 port map ( q=>nx122, i0=>nx3593, i1=>pro_state_11);
   ix113 : an12_x1 port map ( q=>nx112, i0=>nx3591, i1=>pro_state_10);
   ix103 : an12_x1 port map ( q=>nx102, i0=>nx3591, i1=>pro_state_9);
   ix93 : an12_x1 port map ( q=>nx92, i0=>nx3591, i1=>pro_state_8);
   ix83 : an12_x1 port map ( q=>nx82, i0=>nx3591, i1=>pro_state_7);
   ix73 : an12_x1 port map ( q=>nx72, i0=>nx3591, i1=>pro_state_6);
   ix63 : an12_x1 port map ( q=>nx62, i0=>nx3591, i1=>pro_state_5);
   ix53 : an12_x1 port map ( q=>nx52, i0=>nx3589, i1=>pro_state_4);
   ix43 : an12_x1 port map ( q=>nx42, i0=>nx3589, i1=>pro_state_3);
   ix3 : on12_x1 port map ( q=>nx2, i0=>PRO_FUN_parity3_ENABLE, i1=>
      conpro_system_reset);
   ix23 : an12_x1 port map ( q=>nx22, i0=>nx3589, i1=>pro_state_1);
   ix13 : an12_x1 port map ( q=>nx12, i0=>nx3589, i1=>pro_state_0);
   ix709 : o2_x2 port map ( q=>nx708, i0=>pro_state_1, i1=>
      conpro_system_reset);
   ix707 : on12_x4 port map ( q=>nx706, i0=>nx3578, i1=>conpro_system_reset
   );
   ix3588 : on12_x1 port map ( q=>nx3589, i0=>PRO_FUN_parity3_ENABLE, i1=>
      conpro_system_reset);
   ix3590 : on12_x1 port map ( q=>nx3591, i0=>PRO_FUN_parity3_ENABLE, i1=>
      conpro_system_reset);
   ix3592 : on12_x1 port map ( q=>nx3593, i0=>PRO_FUN_parity3_ENABLE, i1=>
      conpro_system_reset);
   ix3594 : on12_x1 port map ( q=>nx3595, i0=>PRO_FUN_parity3_ENABLE, i1=>
      conpro_system_reset);
   ix3596 : on12_x1 port map ( q=>nx3597, i0=>PRO_FUN_parity3_ENABLE, i1=>
      conpro_system_reset);
   ix3598 : on12_x1 port map ( q=>nx3599, i0=>PRO_FUN_parity3_ENABLE, i1=>
      conpro_system_reset);
   ix3600 : on12_x1 port map ( q=>nx3601, i0=>PRO_FUN_parity3_ENABLE, i1=>
      conpro_system_reset);
   ix3602 : on12_x1 port map ( q=>nx3603, i0=>PRO_FUN_parity3_ENABLE, i1=>
      conpro_system_reset);
   ix3604 : on12_x1 port map ( q=>nx3605, i0=>PRO_FUN_parity3_ENABLE, i1=>
      conpro_system_reset);
   ix3606 : on12_x1 port map ( q=>nx3607, i0=>PRO_FUN_parity3_ENABLE, i1=>
      conpro_system_reset);
   ix3608 : on12_x1 port map ( q=>nx3609, i0=>PRO_FUN_parity3_ENABLE, i1=>
      conpro_system_reset);
   ix3618 : o2_x2 port map ( q=>nx3619, i0=>pro_state_1, i1=>
      conpro_system_reset);
   ix3620 : o2_x2 port map ( q=>nx3621, i0=>pro_state_1, i1=>
      conpro_system_reset);
   ix3622 : o2_x2 port map ( q=>nx3623, i0=>pro_state_1, i1=>
      conpro_system_reset);
   ix3624 : o2_x2 port map ( q=>nx3625, i0=>pro_state_1, i1=>
      conpro_system_reset);
   ix3626 : o2_x2 port map ( q=>nx3627, i0=>pro_state_1, i1=>
      conpro_system_reset);
   ix3628 : o2_x2 port map ( q=>nx3629, i0=>pro_state_1, i1=>
      conpro_system_reset);
   ix3630 : o2_x2 port map ( q=>nx3631, i0=>pro_state_1, i1=>
      conpro_system_reset);
   ix3632 : o2_x2 port map ( q=>nx3633, i0=>pro_state_1, i1=>
      conpro_system_reset);
   ix3634 : o2_x2 port map ( q=>nx3635, i0=>pro_state_1, i1=>
      conpro_system_reset);
   ix3636 : o2_x2 port map ( q=>nx3637, i0=>pro_state_1, i1=>
      conpro_system_reset);
   ix3638 : o2_x2 port map ( q=>nx3639, i0=>pro_state_1, i1=>
      conpro_system_reset);
   ix3640 : o2_x2 port map ( q=>nx3641, i0=>pro_state_1, i1=>
      conpro_system_reset);
   ix3642 : o2_x2 port map ( q=>nx3643, i0=>pro_state_1, i1=>
      conpro_system_reset);
   ix3644 : o2_x2 port map ( q=>nx3645, i0=>pro_state_1, i1=>
      conpro_system_reset);
   ix3646 : o2_x2 port map ( q=>nx3647, i0=>pro_state_1, i1=>
      conpro_system_reset);
end main ;

